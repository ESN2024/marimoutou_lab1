
module lab1 (
	clk_clk,
	pio_0_external_connection_export,
	reset_reset_n,
	btn_external_connection_export);	

	input		clk_clk;
	output	[7:0]	pio_0_external_connection_export;
	input		reset_reset_n;
	input		btn_external_connection_export;
endmodule
